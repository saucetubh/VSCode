module priorityencoder_83(input en,input[7:0] inp, output reg[2:0] out);

endmodule