module decoder24_behaviour(input en,input a,input b,output reg[3:0]out);

endmodule