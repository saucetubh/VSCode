module concat;
    wire [3:0] A = 4'b1010;
    wire [3:0] B = 4'b1100; 
    wire [7:0] C;
    
endmodule
