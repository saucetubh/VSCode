module p_encoder(input [3:0]D, output [1:0]Y, output V); //if no input is high, V=0
    
endmodule